module Transform()



endmodule