
module RInitialPermutation(DataIn,DataOut);
	input [63:0] DataIn;
	output [63:0] DataOut;
	assign DataOut[0]=DataIn[39];
	assign DataOut[1]=DataIn[7];
	assign DataOut[2]=DataIn[47];
	assign DataOut[3]=DataIn[15];
	assign DataOut[4]=DataIn[55];
	assign DataOut[5]=DataIn[23];
	assign DataOut[6]=DataIn[63];
	assign DataOut[7]=DataIn[31];
	assign DataOut[8]=DataIn[38];
	assign DataOut[9]=DataIn[6];
	assign DataOut[10]=DataIn[46];
	assign DataOut[11]=DataIn[14];
	assign DataOut[12]=DataIn[54];
	assign DataOut[13]=DataIn[22];
	assign DataOut[14]=DataIn[62];
	assign DataOut[15]=DataIn[30];
	assign DataOut[16]=DataIn[37];
	assign DataOut[17]=DataIn[5];
	assign DataOut[18]=DataIn[45];
	assign DataOut[19]=DataIn[13];
	assign DataOut[20]=DataIn[53];
	assign DataOut[21]=DataIn[21];
	assign DataOut[22]=DataIn[61];
	assign DataOut[23]=DataIn[29];
	assign DataOut[24]=DataIn[36];
	assign DataOut[25]=DataIn[4];
	assign DataOut[26]=DataIn[44];
	assign DataOut[27]=DataIn[12];
	assign DataOut[28]=DataIn[52];
	assign DataOut[29]=DataIn[20];
	assign DataOut[30]=DataIn[60];
	assign DataOut[31]=DataIn[28];
	assign DataOut[32]=DataIn[35];
	assign DataOut[33]=DataIn[3];
	assign DataOut[34]=DataIn[43];
	assign DataOut[35]=DataIn[11];
	assign DataOut[36]=DataIn[51];
	assign DataOut[37]=DataIn[19];
	assign DataOut[38]=DataIn[59];
	assign DataOut[39]=DataIn[27];
	assign DataOut[40]=DataIn[34];
	assign DataOut[41]=DataIn[2];
	assign DataOut[42]=DataIn[42];
	assign DataOut[43]=DataIn[10];
	assign DataOut[44]=DataIn[50];
	assign DataOut[45]=DataIn[18];
	assign DataOut[46]=DataIn[58];
	assign DataOut[47]=DataIn[26];
	assign DataOut[48]=DataIn[33];
	assign DataOut[49]=DataIn[1];
	assign DataOut[50]=DataIn[41];
	assign DataOut[51]=DataIn[9];
	assign DataOut[52]=DataIn[49];
	assign DataOut[53]=DataIn[17];
	assign DataOut[54]=DataIn[57];
	assign DataOut[55]=DataIn[25];
	assign DataOut[56]=DataIn[32];
	assign DataOut[57]=DataIn[0];
	assign DataOut[58]=DataIn[40];
	assign DataOut[59]=DataIn[8];
	assign DataOut[60]=DataIn[48];
	assign DataOut[61]=DataIn[16];
	assign DataOut[62]=DataIn[56];
	assign DataOut[63]=DataIn[24];
endmodule
