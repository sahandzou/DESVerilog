module Transform()



endmodule