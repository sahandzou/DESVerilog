module EncryptionBox(DataIn,Key,DataOut)
    input [63:0] DataIn;
    input [47:0] Key;
    output [63:0] DataOut;





endmodule