module PlainTextitialPermutation(PlaPlainTextText,PermutatedText);
    PlainTextput [63:0] PlaPlainTextText;
    PermutatedTextput [63:0] PermutatedText;
    
    assign PermutatedText[0] = PlainText[57];
    assign PermutatedText[1] = PlainText[49];
    assign PermutatedText[2] = PlainText[41];
    assign PermutatedText[3] = PlainText[33];
    assign PermutatedText[4] = PlainText[25];
    assign PermutatedText[5] = PlainText[17];
    assign PermutatedText[6] = PlainText[9];
    assign PermutatedText[7] = PlainText[1];
    assign PermutatedText[8] = PlainText[59];
    assign PermutatedText[9] = PlainText[51];
    assign PermutatedText[10] = PlainText[43];
    assign PermutatedText[11] = PlainText[35];
    assign PermutatedText[12] = PlainText[27];
    assign PermutatedText[13] = PlainText[19];
    assign PermutatedText[14] = PlainText[11];
    assign PermutatedText[15] = PlainText[3];
    assign PermutatedText[16] = PlainText[61];
    assign PermutatedText[17] = PlainText[53];
    assign PermutatedText[18] = PlainText[45];
    assign PermutatedText[19] = PlainText[37];
    assign PermutatedText[20] = PlainText[29];
    assign PermutatedText[21] = PlainText[21];
    assign PermutatedText[22] = PlainText[13];
    assign PermutatedText[23] = PlainText[5];
    assign PermutatedText[24] = PlainText[63];
    assign PermutatedText[25] = PlainText[55];
    assign PermutatedText[26] = PlainText[47];
    assign PermutatedText[27] = PlainText[39];
    assign PermutatedText[28] = PlainText[31];
    assign PermutatedText[29] = PlainText[23];
    assign PermutatedText[30] = PlainText[15];
    assign PermutatedText[31] = PlainText[7];
    assign PermutatedText[32] = PlainText[56];
    assign PermutatedText[33] = PlainText[48];
    assign PermutatedText[34] = PlainText[40];
    assign PermutatedText[35] = PlainText[32];
    assign PermutatedText[36] = PlainText[24];
    assign PermutatedText[37] = PlainText[16];
    assign PermutatedText[38] = PlainText[8];
    assign PermutatedText[39] = PlainText[0];
    assign PermutatedText[40] = PlainText[58];
    assign PermutatedText[41] = PlainText[50];
    assign PermutatedText[42] = PlainText[42];
    assign PermutatedText[43] = PlainText[34];
    assign PermutatedText[44] = PlainText[26];
    assign PermutatedText[45] = PlainText[18];
    assign PermutatedText[46] = PlainText[10];
    assign PermutatedText[47] = PlainText[2];
    assign PermutatedText[48] = PlainText[60];
    assign PermutatedText[49] = PlainText[52];
    assign PermutatedText[50] = PlainText[44];
    assign PermutatedText[51] = PlainText[36];
    assign PermutatedText[52] = PlainText[28];
    assign PermutatedText[53] = PlainText[20];
    assign PermutatedText[54] = PlainText[12];
    assign PermutatedText[55] = PlainText[4];
    assign PermutatedText[56] = PlainText[62];
    assign PermutatedText[57] = PlainText[54];
    assign PermutatedText[58] = PlainText[46];
    assign PermutatedText[59] = PlainText[38];
    assign PermutatedText[60] = PlainText[30];
    assign PermutatedText[61] = PlainText[22];
    assign PermutatedText[62] = PlainText[14];
    assign PermutatedText[63] = PlainText[9];

endmoudle